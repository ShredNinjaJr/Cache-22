package L1_cache_types;

typedef logic [8:0] cache_tag;
typedef logic [2:0] cache_index;
typedef logic [2:0] cache_offset;

endpackage
