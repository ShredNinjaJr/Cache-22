import lc3b_types::*;

module mp3
(
	input clk
);


 
 endmodule: mp3